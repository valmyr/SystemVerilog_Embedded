module adpcm()

endmodule
